module counter #(
    
) (
    input wire pulse_1,
    input wire pulse_2,
    input wire pulse_3,
    input wire clk,
    output reg [16]counter

);

always @(posedge clk) begin
    
end

endmodule
